test hoi
